`define flit_size 32
`define router_address_size 5
`define flit_num_beg_index 
`define flit_num_end_index
`define address_beg_index
`define address_end_index
`define type_beg_index
`define type_end_index


module utils ;
  