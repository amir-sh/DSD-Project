`define flit_size 32
`define router_address_size 5
`define flit_num_beg_index 
`define flit_num_end_index
`define package_size_beg_index 24 
`define package_size_end_index 22
`define dest_address_beg_index
`define dest_address_end_index
`define type_beg_index
`define type_end_index


module utils ;
  